`timescale 1ns / 10ps

module signed_multiplier #(
    // parameters
) (
    input clk, n_rst
);



endmodule


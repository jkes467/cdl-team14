`timescale 1ns / 10ps

module multiply_by_2 #(
    // parameters
) (
    input clk, n_rst
);



endmodule


`timescale 1ns / 10ps

module controller #(
    // parameters
) (
    input clk, n_rst
);



endmodule


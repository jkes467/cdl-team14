`timescale 1ns / 10ps

module ai_accelerator #(
    // parameters
) (
    input clk, n_rst
);



endmodule


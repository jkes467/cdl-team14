`timescale 1ns / 10ps

module sram_buffer #(
    // parameters
) (
    input clk, n_rst
);



endmodule


`timescale 1ns / 10ps

module systolic_array #(
    // parameters
) (
    input clk, n_rst
);



endmodule


`timescale 1ns / 10ps

module PE #(
    // parameters
) (
    input clk, n_rst
);



endmodule


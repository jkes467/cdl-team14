`timescale 1ns / 10ps

module bias_adder #(
    // parameters
) (
    input clk, n_rst
);



endmodule


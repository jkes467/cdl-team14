`timescale 1ns / 10ps

module activation #(
    // parameters
) (
    input clk, n_rst
);



endmodule

